module top_module(Hclk,Hresetn,Hwrite,Hreadyin,Hreadyout,Hwdata,Haddr,Htrans,Prdata,Penable,Pwrite,Pselx,Paddr,Pwdata,Hreadyout,Hresp,Hrdata);

 input Hclk,Hresetn,Hwrite,Hreadyin;
 input [31:0] Hwdata,Haddr,Prdata;
 input[1:0] Htrans;
 output Penable,Pwrite,Hreadyout;
 output [1:0] Hresp; 
 output [2:0] Pselx;
 output [31:0] Paddr,Pwdata;
 output [31:0] Hrdata;

///////////////////////////////////////////////////////////////INTERMEDIATE SIGNALS

 wire valid;
 wire [31:0] Haddr1,Haddr2,Hwdata1,Hwdata2;
 wire Hwritereg;
 wire [2:0] tempselx;

/////////////////////////////////////////////////////////////// MODULE INSTANTIATIONS


 ahb_slave_interface apbslave (Hclk,Hresetn,Hwrite,Hreadyin,Htrans,Haddr,Hwdata,Prdata,valid,Haddr1,Haddr2,Hwdata1,Hwdata2,Hrdata,Hwritereg,tempselx,Hresp);


 apb_fsm_controller apbcontrol (Hclk,Hresetn,valid,Haddr1,Haddr2,Hwdata1,Hwdata2,Prdata,Hwrite,Haddr,Hwdata,Hwritereg,tempselx,Pwrite,Penable,Pselx,Paddr,Pwdata,Hreadyout);


endmodule

